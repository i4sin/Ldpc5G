package BASE_TEST;
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    `include "BaseTest.svh"
endpackage
