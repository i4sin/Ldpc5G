package SEQUENCE;
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    `include "Seq.svh"
endpackage
