module LdpcLoopWrapper (
    AxisIf.slave s_axis,
    AxisIf.master m_axis
);
    
endmodule
