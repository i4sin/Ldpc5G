package RANGE;
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    `include "Range.svh"
endpackage
