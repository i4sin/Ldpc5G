package AXIS_CONNECTOR_TEST;
    import vunit_pkg::*;
    `include "vunit_defines.svh"

    `include "Env.svh"
endpackage
