package TEST_CASES;
    import uvm_pkg::*;
    `include "uvm_macros.svh"
    
    import AXIS_CONNECTOR_TEST::*;
    import AXIS_VIP::*;
    import BASE_TEST::*;
    import CONFIG_DB::*;
    import RESET_VIP::*;

    `include "Test.svh"
endpackage
