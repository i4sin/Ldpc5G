package ANALYSIS_MAP;
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    `include "AnalysisMap.svh"
    `include "AnalysisCastMap.svh"
endpackage
