interface ClockIf (
    input clk
);
endinterface
