interface ClockIf;
    logic clk;
endinterface
