package TEST_CASES;
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    `include "Test.svh"
endpackage
