package DRIVER;
    import uvm_pkg::*;
    `include "uvm_macros.svh"
    
    import CONFIG_DB::*;

    `include "Driver.svh"
endpackage
