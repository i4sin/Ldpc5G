interface ResetIf (
    input aclk
);
    logic aresetn;
endinterface
