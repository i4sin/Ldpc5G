package CONFIG_DB;
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    `include "ConfigDb.svh"
endpackage