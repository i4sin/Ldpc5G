package WATCHDOG;
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    `include "Watchdog.svh"
endpackage
