package RESET_VIP;
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    `include "ResetItem.svh"
    `include "ResetPacket.svh"
    `include "InitialResetSeq.svh"
    
    `include "ResetDriver.svh"
    `include "ResetSeqr.svh"
    `include "ResetAgent.svh"
endpackage
