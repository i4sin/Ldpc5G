package SEQUENCE;
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    import CONFIG_DB::*;

    `include "Item.svh"
    `include "Seq.svh"
    `include "RepeatSeq.svh"
    `include "CountSeq.svh"
    `include "InfiniteSeq.svh"
endpackage
