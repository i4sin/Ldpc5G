package AXIS_VIP;
    import uvm::*;
    `include "uvm_macros.svh"

    `include "AxisMasterItem.svh"
    `include "AxisMasterPacket.svh"
    `include "AxisTransaction.svh"
    
    `include "AxisMasterDriver.svh"
    `include "AxisMonitor.svh"
endpackage