package TEST_CASES;
    import vunit_pkg::*;
    `include "vunit_defines.svh"

    `include "Test.svh"
endpackage
