package BASE_TEST;
    import uvm_pkg::*;
    `include "uvm_macros.svh"
    
    import CONFIG_DB::*;
    import WATCHDOG::*;

    `include "BaseTest.svh"
endpackage
