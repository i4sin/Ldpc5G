package LDPC_LOOP_WRAPPER_TEST;
    import uvm_pkg::*;
    `include "uvm_macros.svh"
    
    import AXIS_VIP::*;
    import CONFIG_DB::*;
    import RESET_VIP::*;

    `include "ControlCfg.svh"

    `include "DecoderControlItem.svh"
    `include "EncoderControlItem.svh"

    `include "Scoreboard.svh"
    `include "Env.svh"
endpackage
