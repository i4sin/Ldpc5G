package AXIS_CONNECTOR_TEST;
    import uvm_pkg::*;
    `include "uvm_macros.svh"
    
    import AXIS_VIP::*;
    import CONFIG_DB::*;
    import RESET_VIP::*;

    `include "Scoreboard.svh"
    `include "Env.svh"
endpackage
