package AXIS_CONNECTOR_TEST;
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    `include "Env.svh"
    `include "Scoreboard.svh"
endpackage
