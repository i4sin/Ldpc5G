interface ResetIf (
    input clk
);
    logic resetn;
endinterface
