package LDPC_LOOP_WRAPPER_TEST;
    import uvm_pkg::*;
    `include "uvm_macros.svh"
    
    import AXIS_VIP::*;
    import CONFIG_DB::*;
    import LDPC_IP_CONTROL_PKG::*;
    import RESET_VIP::*;

    `include "AxisMasterDecoderControlItem.svh"
    `include "AxisMasterEncoderControlItem.svh"

    `include "Scoreboard.svh"
    `include "Env.svh"
endpackage
