package MONITOR;
    import uvm_pkg::*;
    `include "uvm_macros.svh"
    
    import CONFIG_DB::*;

    `include "Monitor.svh"
endpackage
