package WATCHDOG;
    import uvm_pkg::*;
    `include "uvm_macros.svh"
    
    import CONFIG_DB::*;

    `include "Watchdog.svh"
endpackage
