package RESET_VIP;
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    import CONFIG_DB::*;
    import SEQUENCE::*;

    `include "ResetItem.svh"
    `include "InitialResetSeq.svh"
    
    `include "ResetDriver.svh"
    `include "ResetSeqr.svh"
    `include "ResetAgent.svh"
endpackage
