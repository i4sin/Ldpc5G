package AXIS_VIP;
    import uvm::*;
    `include "uvm_macros.svh"

    `include "AxisMasterItem.svh"
    `include "AxisMasterPacket.svh"
    `include "AxisMasterPacketSeq.svh"
    `include "AxisTransaction.svh"
    
    `include "AxisMasterDriver.svh"
    `include "AxisMasterSequencer.svh"
    `include "AxisMonitor.svh"
endpackage